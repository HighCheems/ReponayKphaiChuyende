
module CONV_2D_4_Kernel_3_Channel_7 #(
parameter IMG_Width=7, 
parameter IMG_Height=7, 
parameter Datawidth=16, 
parameter Stride=2,
parameter ReLU=1,
parameter w000 = 1,
parameter w010 = 1,
parameter w020 = 1,
parameter w001 = 1,
parameter w011 = 1,
parameter w021 = 1,
parameter w002 = 1,
parameter w012 = 1,
parameter w022 = 1,
parameter w003 = 1,
parameter w013 = 1,
parameter w023 = 1,
parameter w004 = 1,
parameter w014 = 1,
parameter w024 = 1,
parameter w005 = 1,
parameter w015 = 1,
parameter w025 = 1,
parameter w006 = 1,
parameter w016 = 1,
parameter w026 = 1,
parameter w007 = 1,
parameter w017 = 1,
parameter w027 = 1,
parameter w008 = 1,
parameter w018 = 1,
parameter w028 = 1,
parameter w009 = 1,
parameter w019 = 1,
parameter w029 = 1,
parameter w0010 = 1,
parameter w0110 = 1,
parameter w0210 = 1,
parameter w0011 = 1,
parameter w0111 = 1,
parameter w0211 = 1,
parameter w0012 = 1,
parameter w0112 = 1,
parameter w0212 = 1,
parameter w0013 = 1,
parameter w0113 = 1,
parameter w0213 = 1,
parameter w0014 = 1,
parameter w0114 = 1,
parameter w0214 = 1,
parameter w0015 = 1,
parameter w0115 = 1,
parameter w0215 = 1,
parameter w0016 = 1,
parameter w0116 = 1,
parameter w0216 = 1,
parameter w0017 = 1,
parameter w0117 = 1,
parameter w0217 = 1,
parameter w0018 = 1,
parameter w0118 = 1,
parameter w0218 = 1,
parameter w0019 = 1,
parameter w0119 = 1,
parameter w0219 = 1,
parameter w0020 = 1,
parameter w0120 = 1,
parameter w0220 = 1,
parameter w0021 = 1,
parameter w0121 = 1,
parameter w0221 = 1,
parameter w0022 = 1,
parameter w0122 = 1,
parameter w0222 = 1,
parameter w0023 = 1,
parameter w0123 = 1,
parameter w0223 = 1,
parameter w0024 = 1,
parameter w0124 = 1,
parameter w0224 = 1,
parameter w0025 = 1,
parameter w0125 = 1,
parameter w0225 = 1,
parameter w0026 = 1,
parameter w0126 = 1,
parameter w0226 = 1,
parameter w0027 = 1,
parameter w0127 = 1,
parameter w0227 = 1,
parameter w0028 = 1,
parameter w0128 = 1,
parameter w0228 = 1,
parameter w0029 = 1,
parameter w0129 = 1,
parameter w0229 = 1,
parameter w0030 = 1,
parameter w0130 = 1,
parameter w0230 = 1,
parameter w0031 = 1,
parameter w0131 = 1,
parameter w0231 = 1,
parameter w0032 = 1,
parameter w0132 = 1,
parameter w0232 = 1,
parameter w0033 = 1,
parameter w0133 = 1,
parameter w0233 = 1,
parameter w0034 = 1,
parameter w0134 = 1,
parameter w0234 = 1,
parameter w0035 = 1,
parameter w0135 = 1,
parameter w0235 = 1,
parameter w0036 = 1,
parameter w0136 = 1,
parameter w0236 = 1,
parameter w0037 = 1,
parameter w0137 = 1,
parameter w0237 = 1,
parameter w0038 = 1,
parameter w0138 = 1,
parameter w0238 = 1,
parameter w0039 = 1,
parameter w0139 = 1,
parameter w0239 = 1,
parameter w0040 = 1,
parameter w0140 = 1,
parameter w0240 = 1,
parameter w0041 = 1,
parameter w0141 = 1,
parameter w0241 = 1,
parameter w0042 = 1,
parameter w0142 = 1,
parameter w0242 = 1,
parameter w0043 = 1,
parameter w0143 = 1,
parameter w0243 = 1,
parameter w0044 = 1,
parameter w0144 = 1,
parameter w0244 = 1,
parameter w0045 = 1,
parameter w0145 = 1,
parameter w0245 = 1,
parameter w0046 = 1,
parameter w0146 = 1,
parameter w0246 = 1,
parameter w0047 = 1,
parameter w0147 = 1,
parameter w0247 = 1,
parameter w0048 = 1,
parameter w0148 = 1,
parameter w0248 = 1,
parameter bias_0 = 1,
parameter w100 = 1,
parameter w110 = 1,
parameter w120 = 1,
parameter w101 = 1,
parameter w111 = 1,
parameter w121 = 1,
parameter w102 = 1,
parameter w112 = 1,
parameter w122 = 1,
parameter w103 = 1,
parameter w113 = 1,
parameter w123 = 1,
parameter w104 = 1,
parameter w114 = 1,
parameter w124 = 1,
parameter w105 = 1,
parameter w115 = 1,
parameter w125 = 1,
parameter w106 = 1,
parameter w116 = 1,
parameter w126 = 1,
parameter w107 = 1,
parameter w117 = 1,
parameter w127 = 1,
parameter w108 = 1,
parameter w118 = 1,
parameter w128 = 1,
parameter w109 = 1,
parameter w119 = 1,
parameter w129 = 1,
parameter w1010 = 1,
parameter w1110 = 1,
parameter w1210 = 1,
parameter w1011 = 1,
parameter w1111 = 1,
parameter w1211 = 1,
parameter w1012 = 1,
parameter w1112 = 1,
parameter w1212 = 1,
parameter w1013 = 1,
parameter w1113 = 1,
parameter w1213 = 1,
parameter w1014 = 1,
parameter w1114 = 1,
parameter w1214 = 1,
parameter w1015 = 1,
parameter w1115 = 1,
parameter w1215 = 1,
parameter w1016 = 1,
parameter w1116 = 1,
parameter w1216 = 1,
parameter w1017 = 1,
parameter w1117 = 1,
parameter w1217 = 1,
parameter w1018 = 1,
parameter w1118 = 1,
parameter w1218 = 1,
parameter w1019 = 1,
parameter w1119 = 1,
parameter w1219 = 1,
parameter w1020 = 1,
parameter w1120 = 1,
parameter w1220 = 1,
parameter w1021 = 1,
parameter w1121 = 1,
parameter w1221 = 1,
parameter w1022 = 1,
parameter w1122 = 1,
parameter w1222 = 1,
parameter w1023 = 1,
parameter w1123 = 1,
parameter w1223 = 1,
parameter w1024 = 1,
parameter w1124 = 1,
parameter w1224 = 1,
parameter w1025 = 1,
parameter w1125 = 1,
parameter w1225 = 1,
parameter w1026 = 1,
parameter w1126 = 1,
parameter w1226 = 1,
parameter w1027 = 1,
parameter w1127 = 1,
parameter w1227 = 1,
parameter w1028 = 1,
parameter w1128 = 1,
parameter w1228 = 1,
parameter w1029 = 1,
parameter w1129 = 1,
parameter w1229 = 1,
parameter w1030 = 1,
parameter w1130 = 1,
parameter w1230 = 1,
parameter w1031 = 1,
parameter w1131 = 1,
parameter w1231 = 1,
parameter w1032 = 1,
parameter w1132 = 1,
parameter w1232 = 1,
parameter w1033 = 1,
parameter w1133 = 1,
parameter w1233 = 1,
parameter w1034 = 1,
parameter w1134 = 1,
parameter w1234 = 1,
parameter w1035 = 1,
parameter w1135 = 1,
parameter w1235 = 1,
parameter w1036 = 1,
parameter w1136 = 1,
parameter w1236 = 1,
parameter w1037 = 1,
parameter w1137 = 1,
parameter w1237 = 1,
parameter w1038 = 1,
parameter w1138 = 1,
parameter w1238 = 1,
parameter w1039 = 1,
parameter w1139 = 1,
parameter w1239 = 1,
parameter w1040 = 1,
parameter w1140 = 1,
parameter w1240 = 1,
parameter w1041 = 1,
parameter w1141 = 1,
parameter w1241 = 1,
parameter w1042 = 1,
parameter w1142 = 1,
parameter w1242 = 1,
parameter w1043 = 1,
parameter w1143 = 1,
parameter w1243 = 1,
parameter w1044 = 1,
parameter w1144 = 1,
parameter w1244 = 1,
parameter w1045 = 1,
parameter w1145 = 1,
parameter w1245 = 1,
parameter w1046 = 1,
parameter w1146 = 1,
parameter w1246 = 1,
parameter w1047 = 1,
parameter w1147 = 1,
parameter w1247 = 1,
parameter w1048 = 1,
parameter w1148 = 1,
parameter w1248 = 1,
parameter bias_1 = 2,
parameter w200 = 1,
parameter w210 = 1,
parameter w220 = 1,
parameter w201 = 1,
parameter w211 = 1,
parameter w221 = 1,
parameter w202 = 1,
parameter w212 = 1,
parameter w222 = 1,
parameter w203 = 1,
parameter w213 = 1,
parameter w223 = 1,
parameter w204 = 1,
parameter w214 = 1,
parameter w224 = 1,
parameter w205 = 1,
parameter w215 = 1,
parameter w225 = 1,
parameter w206 = 1,
parameter w216 = 1,
parameter w226 = 1,
parameter w207 = 1,
parameter w217 = 1,
parameter w227 = 1,
parameter w208 = 1,
parameter w218 = 1,
parameter w228 = 1,
parameter w209 = 1,
parameter w219 = 1,
parameter w229 = 1,
parameter w2010 = 1,
parameter w2110 = 1,
parameter w2210 = 1,
parameter w2011 = 1,
parameter w2111 = 1,
parameter w2211 = 1,
parameter w2012 = 1,
parameter w2112 = 1,
parameter w2212 = 1,
parameter w2013 = 1,
parameter w2113 = 1,
parameter w2213 = 1,
parameter w2014 = 1,
parameter w2114 = 1,
parameter w2214 = 1,
parameter w2015 = 1,
parameter w2115 = 1,
parameter w2215 = 1,
parameter w2016 = 1,
parameter w2116 = 1,
parameter w2216 = 1,
parameter w2017 = 1,
parameter w2117 = 1,
parameter w2217 = 1,
parameter w2018 = 1,
parameter w2118 = 1,
parameter w2218 = 1,
parameter w2019 = 1,
parameter w2119 = 1,
parameter w2219 = 1,
parameter w2020 = 1,
parameter w2120 = 1,
parameter w2220 = 1,
parameter w2021 = 1,
parameter w2121 = 1,
parameter w2221 = 1,
parameter w2022 = 1,
parameter w2122 = 1,
parameter w2222 = 1,
parameter w2023 = 1,
parameter w2123 = 1,
parameter w2223 = 1,
parameter w2024 = 1,
parameter w2124 = 1,
parameter w2224 = 1,
parameter w2025 = 1,
parameter w2125 = 1,
parameter w2225 = 1,
parameter w2026 = 1,
parameter w2126 = 1,
parameter w2226 = 1,
parameter w2027 = 1,
parameter w2127 = 1,
parameter w2227 = 1,
parameter w2028 = 1,
parameter w2128 = 1,
parameter w2228 = 1,
parameter w2029 = 1,
parameter w2129 = 1,
parameter w2229 = 1,
parameter w2030 = 1,
parameter w2130 = 1,
parameter w2230 = 1,
parameter w2031 = 1,
parameter w2131 = 1,
parameter w2231 = 1,
parameter w2032 = 1,
parameter w2132 = 1,
parameter w2232 = 1,
parameter w2033 = 1,
parameter w2133 = 1,
parameter w2233 = 1,
parameter w2034 = 1,
parameter w2134 = 1,
parameter w2234 = 1,
parameter w2035 = 1,
parameter w2135 = 1,
parameter w2235 = 1,
parameter w2036 = 1,
parameter w2136 = 1,
parameter w2236 = 1,
parameter w2037 = 1,
parameter w2137 = 1,
parameter w2237 = 1,
parameter w2038 = 1,
parameter w2138 = 1,
parameter w2238 = 1,
parameter w2039 = 1,
parameter w2139 = 1,
parameter w2239 = 1,
parameter w2040 = 1,
parameter w2140 = 1,
parameter w2240 = 1,
parameter w2041 = 1,
parameter w2141 = 1,
parameter w2241 = 1,
parameter w2042 = 1,
parameter w2142 = 1,
parameter w2242 = 1,
parameter w2043 = 1,
parameter w2143 = 1,
parameter w2243 = 1,
parameter w2044 = 1,
parameter w2144 = 1,
parameter w2244 = 1,
parameter w2045 = 1,
parameter w2145 = 1,
parameter w2245 = 1,
parameter w2046 = 1,
parameter w2146 = 1,
parameter w2246 = 1,
parameter w2047 = 1,
parameter w2147 = 1,
parameter w2247 = 1,
parameter w2048 = 1,
parameter w2148 = 1,
parameter w2248 = 1,
parameter bias_2 = 3,
parameter w300 = 1,
parameter w310 = 1,
parameter w320 = 1,
parameter w301 = 1,
parameter w311 = 1,
parameter w321 = 1,
parameter w302 = 1,
parameter w312 = 1,
parameter w322 = 1,
parameter w303 = 1,
parameter w313 = 1,
parameter w323 = 1,
parameter w304 = 1,
parameter w314 = 1,
parameter w324 = 1,
parameter w305 = 1,
parameter w315 = 1,
parameter w325 = 1,
parameter w306 = 1,
parameter w316 = 1,
parameter w326 = 1,
parameter w307 = 1,
parameter w317 = 1,
parameter w327 = 1,
parameter w308 = 1,
parameter w318 = 1,
parameter w328 = 1,
parameter w309 = 1,
parameter w319 = 1,
parameter w329 = 1,
parameter w3010 = 1,
parameter w3110 = 1,
parameter w3210 = 1,
parameter w3011 = 1,
parameter w3111 = 1,
parameter w3211 = 1,
parameter w3012 = 1,
parameter w3112 = 1,
parameter w3212 = 1,
parameter w3013 = 1,
parameter w3113 = 1,
parameter w3213 = 1,
parameter w3014 = 1,
parameter w3114 = 1,
parameter w3214 = 1,
parameter w3015 = 1,
parameter w3115 = 1,
parameter w3215 = 1,
parameter w3016 = 1,
parameter w3116 = 1,
parameter w3216 = 1,
parameter w3017 = 1,
parameter w3117 = 1,
parameter w3217 = 1,
parameter w3018 = 1,
parameter w3118 = 1,
parameter w3218 = 1,
parameter w3019 = 1,
parameter w3119 = 1,
parameter w3219 = 1,
parameter w3020 = 1,
parameter w3120 = 1,
parameter w3220 = 1,
parameter w3021 = 1,
parameter w3121 = 1,
parameter w3221 = 1,
parameter w3022 = 1,
parameter w3122 = 1,
parameter w3222 = 1,
parameter w3023 = 1,
parameter w3123 = 1,
parameter w3223 = 1,
parameter w3024 = 1,
parameter w3124 = 1,
parameter w3224 = 1,
parameter w3025 = 1,
parameter w3125 = 1,
parameter w3225 = 1,
parameter w3026 = 1,
parameter w3126 = 1,
parameter w3226 = 1,
parameter w3027 = 1,
parameter w3127 = 1,
parameter w3227 = 1,
parameter w3028 = 1,
parameter w3128 = 1,
parameter w3228 = 1,
parameter w3029 = 1,
parameter w3129 = 1,
parameter w3229 = 1,
parameter w3030 = 1,
parameter w3130 = 1,
parameter w3230 = 1,
parameter w3031 = 1,
parameter w3131 = 1,
parameter w3231 = 1,
parameter w3032 = 1,
parameter w3132 = 1,
parameter w3232 = 1,
parameter w3033 = 1,
parameter w3133 = 1,
parameter w3233 = 1,
parameter w3034 = 1,
parameter w3134 = 1,
parameter w3234 = 1,
parameter w3035 = 1,
parameter w3135 = 1,
parameter w3235 = 1,
parameter w3036 = 1,
parameter w3136 = 1,
parameter w3236 = 1,
parameter w3037 = 1,
parameter w3137 = 1,
parameter w3237 = 1,
parameter w3038 = 1,
parameter w3138 = 1,
parameter w3238 = 1,
parameter w3039 = 1,
parameter w3139 = 1,
parameter w3239 = 1,
parameter w3040 = 1,
parameter w3140 = 1,
parameter w3240 = 1,
parameter w3041 = 1,
parameter w3141 = 1,
parameter w3241 = 1,
parameter w3042 = 1,
parameter w3142 = 1,
parameter w3242 = 1,
parameter w3043 = 1,
parameter w3143 = 1,
parameter w3243 = 1,
parameter w3044 = 1,
parameter w3144 = 1,
parameter w3244 = 1,
parameter w3045 = 1,
parameter w3145 = 1,
parameter w3245 = 1,
parameter w3046 = 1,
parameter w3146 = 1,
parameter w3246 = 1,
parameter w3047 = 1,
parameter w3147 = 1,
parameter w3247 = 1,
parameter w3048 = 1,
parameter w3148 = 1,
parameter w3248 = 1,
parameter bias_3 = 4

)
(
clk,rst,valid_in,
In_0,
In_1,
In_2,
valid_out,
Out_0,
Out_1,
Out_2,
Out_3
);

// port map
input wire clk,rst,valid_in;
input wire [Datawidth-1:0] In_0,In_1,In_2;
output reg valid_out;
output reg [Datawidth-1:0] Out_0;
output reg [Datawidth-1:0] Out_1;
output reg [Datawidth-1:0] Out_2;
output reg [Datawidth-1:0] Out_3;

wire [Datawidth-1:0] save_Out_0,save_Out_1,save_Out_2,save_Out_3;
wire valid_out_0,valid_out_1,valid_out_2,valid_out_3;
// clk
always @(posedge clk) begin
	if(rst==1'd1) begin
		valid_out<=1'd0;
		Out_0<={Datawidth{1'b0}};
		Out_1<={Datawidth{1'b0}};	
		Out_2<={Datawidth{1'b0}};
		Out_3<={Datawidth{1'b0}};
	end
	else begin
		if(valid_out_0 ==1'd1 && valid_out_1 ==1'd1 && valid_out_2 ==1'd1 && valid_out_3 ==1'd1) begin
			Out_0<=save_Out_0;
			Out_1<=save_Out_1;	
			Out_2<=save_Out_2;
			Out_3<=save_Out_3;
			valid_out<=1'd1;
		end
		else begin
		valid_out<=1'd0;
		end
	end
end

 
CONV_2D_1_Kernel_3_Channel_7 #(
.IMG_Width(IMG_Width), 
.IMG_Height(IMG_Height), 
.Datawidth(Datawidth), 
.Stride(Stride),
.ReLU(ReLU),
.w00(w000),
.w01(w001),
.w02(w002),
.w03(w003),
.w04(w004),
.w05(w005),
.w06(w006),
.w07(w007),
.w08(w008),
.w09(w009),
.w010(w0010),
.w011(w0011),
.w012(w0012),
.w013(w0013),
.w014(w0014),
.w015(w0015),
.w016(w0016),
.w017(w0017),
.w018(w0018),
.w019(w0019),
.w020(w0020),
.w021(w0021),
.w022(w0022),
.w023(w0023),
.w024(w0024),
.w025(w0025),
.w026(w0026),
.w027(w0027),
.w028(w0028),
.w029(w0029),
.w030(w0030),
.w031(w0031),
.w032(w0032),
.w033(w0033),
.w034(w0034),
.w035(w0035),
.w036(w0036),
.w037(w0037),
.w038(w0038),
.w039(w0039),
.w040(w0040),
.w041(w0041),
.w042(w0042),
.w043(w0043),
.w044(w0044),
.w045(w0045),
.w046(w0046),
.w047(w0047),
.w048(w0048),
.w10(w010),
.w11(w011),
.w12(w012),
.w13(w013),
.w14(w014),
.w15(w015),
.w16(w016),
.w17(w017),
.w18(w018),
.w19(w019),
.w110(w0110),
.w111(w0111),
.w112(w0112),
.w113(w0113),
.w114(w0114),
.w115(w0115),
.w116(w0116),
.w117(w0117),
.w118(w0118),
.w119(w0119),
.w120(w0120),
.w121(w0121),
.w122(w0122),
.w123(w0123),
.w124(w0124),
.w125(w0125),
.w126(w0126),
.w127(w0127),
.w128(w0128),
.w129(w0129),
.w130(w0130),
.w131(w0131),
.w132(w0132),
.w133(w0133),
.w134(w0134),
.w135(w0135),
.w136(w0136),
.w137(w0137),
.w138(w0138),
.w139(w0139),
.w140(w0140),
.w141(w0141),
.w142(w0142),
.w143(w0143),
.w144(w0144),
.w145(w0145),
.w146(w0146),
.w147(w0147),
.w148(w0148),
.w20(w020),
.w21(w021),
.w22(w022),
.w23(w023),
.w24(w024),
.w25(w025),
.w26(w026),
.w27(w027),
.w28(w028),
.w29(w029),
.w210(w0210),
.w211(w0211),
.w212(w0212),
.w213(w0213),
.w214(w0214),
.w215(w0215),
.w216(w0216),
.w217(w0217),
.w218(w0218),
.w219(w0219),
.w220(w0220),
.w221(w0221),
.w222(w0222),
.w223(w0223),
.w224(w0224),
.w225(w0225),
.w226(w0226),
.w227(w0227),
.w228(w0228),
.w229(w0229),
.w230(w0230),
.w231(w0231),
.w232(w0232),
.w233(w0233),
.w234(w0234),
.w235(w0235),
.w236(w0236),
.w237(w0237),
.w238(w0238),
.w239(w0239),
.w240(w0240),
.w241(w0241),
.w242(w0242),
.w243(w0243),
.w244(w0244),
.w245(w0245),
.w246(w0246),
.w247(w0247),
.w248(w0248),
.bias(bias_0)
) block_1kernel_0
(
.clk(clk),
.rst(rst),
.valid_in(valid_in),
.In_0(In_0),
.In_1(In_1),
.In_2(In_2),
.Out(save_Out_0),
.valid_out(valid_out_0)
);

 
CONV_2D_1_Kernel_3_Channel_7 #(
.IMG_Width(IMG_Width), 
.IMG_Height(IMG_Height), 
.Datawidth(Datawidth), 
.Stride(Stride),
.ReLU(ReLU),
.w00(w100),
.w01(w101),
.w02(w102),
.w03(w103),
.w04(w104),
.w05(w105),
.w06(w106),
.w07(w107),
.w08(w108),
.w09(w109),
.w010(w1010),
.w011(w1011),
.w012(w1012),
.w013(w1013),
.w014(w1014),
.w015(w1015),
.w016(w1016),
.w017(w1017),
.w018(w1018),
.w019(w1019),
.w020(w1020),
.w021(w1021),
.w022(w1022),
.w023(w1023),
.w024(w1024),
.w025(w1025),
.w026(w1026),
.w027(w1027),
.w028(w1028),
.w029(w1029),
.w030(w1030),
.w031(w1031),
.w032(w1032),
.w033(w1033),
.w034(w1034),
.w035(w1035),
.w036(w1036),
.w037(w1037),
.w038(w1038),
.w039(w1039),
.w040(w1040),
.w041(w1041),
.w042(w1042),
.w043(w1043),
.w044(w1044),
.w045(w1045),
.w046(w1046),
.w047(w1047),
.w048(w1048),
.w10(w110),
.w11(w111),
.w12(w112),
.w13(w113),
.w14(w114),
.w15(w115),
.w16(w116),
.w17(w117),
.w18(w118),
.w19(w119),
.w110(w1110),
.w111(w1111),
.w112(w1112),
.w113(w1113),
.w114(w1114),
.w115(w1115),
.w116(w1116),
.w117(w1117),
.w118(w1118),
.w119(w1119),
.w120(w1120),
.w121(w1121),
.w122(w1122),
.w123(w1123),
.w124(w1124),
.w125(w1125),
.w126(w1126),
.w127(w1127),
.w128(w1128),
.w129(w1129),
.w130(w1130),
.w131(w1131),
.w132(w1132),
.w133(w1133),
.w134(w1134),
.w135(w1135),
.w136(w1136),
.w137(w1137),
.w138(w1138),
.w139(w1139),
.w140(w1140),
.w141(w1141),
.w142(w1142),
.w143(w1143),
.w144(w1144),
.w145(w1145),
.w146(w1146),
.w147(w1147),
.w148(w1148),
.w20(w120),
.w21(w121),
.w22(w122),
.w23(w123),
.w24(w124),
.w25(w125),
.w26(w126),
.w27(w127),
.w28(w128),
.w29(w129),
.w210(w1210),
.w211(w1211),
.w212(w1212),
.w213(w1213),
.w214(w1214),
.w215(w1215),
.w216(w1216),
.w217(w1217),
.w218(w1218),
.w219(w1219),
.w220(w1220),
.w221(w1221),
.w222(w1222),
.w223(w1223),
.w224(w1224),
.w225(w1225),
.w226(w1226),
.w227(w1227),
.w228(w1228),
.w229(w1229),
.w230(w1230),
.w231(w1231),
.w232(w1232),
.w233(w1233),
.w234(w1234),
.w235(w1235),
.w236(w1236),
.w237(w1237),
.w238(w1238),
.w239(w1239),
.w240(w1240),
.w241(w1241),
.w242(w1242),
.w243(w1243),
.w244(w1244),
.w245(w1245),
.w246(w1246),
.w247(w1247),
.w248(w1248),
.bias(bias_1)
) block_1kernel_1
(
.clk(clk),
.rst(rst),
.valid_in(valid_in),
.In_0(In_0),
.In_1(In_1),
.In_2(In_2),
.Out(save_Out_1),
.valid_out(valid_out_1)
);

 
CONV_2D_1_Kernel_3_Channel_7 #(
.IMG_Width(IMG_Width), 
.IMG_Height(IMG_Height), 
.Datawidth(Datawidth), 
.Stride(Stride),
.ReLU(ReLU),
.w00(w200),
.w01(w201),
.w02(w202),
.w03(w203),
.w04(w204),
.w05(w205),
.w06(w206),
.w07(w207),
.w08(w208),
.w09(w209),
.w010(w2010),
.w011(w2011),
.w012(w2012),
.w013(w2013),
.w014(w2014),
.w015(w2015),
.w016(w2016),
.w017(w2017),
.w018(w2018),
.w019(w2019),
.w020(w2020),
.w021(w2021),
.w022(w2022),
.w023(w2023),
.w024(w2024),
.w025(w2025),
.w026(w2026),
.w027(w2027),
.w028(w2028),
.w029(w2029),
.w030(w2030),
.w031(w2031),
.w032(w2032),
.w033(w2033),
.w034(w2034),
.w035(w2035),
.w036(w2036),
.w037(w2037),
.w038(w2038),
.w039(w2039),
.w040(w2040),
.w041(w2041),
.w042(w2042),
.w043(w2043),
.w044(w2044),
.w045(w2045),
.w046(w2046),
.w047(w2047),
.w048(w2048),
.w10(w210),
.w11(w211),
.w12(w212),
.w13(w213),
.w14(w214),
.w15(w215),
.w16(w216),
.w17(w217),
.w18(w218),
.w19(w219),
.w110(w2110),
.w111(w2111),
.w112(w2112),
.w113(w2113),
.w114(w2114),
.w115(w2115),
.w116(w2116),
.w117(w2117),
.w118(w2118),
.w119(w2119),
.w120(w2120),
.w121(w2121),
.w122(w2122),
.w123(w2123),
.w124(w2124),
.w125(w2125),
.w126(w2126),
.w127(w2127),
.w128(w2128),
.w129(w2129),
.w130(w2130),
.w131(w2131),
.w132(w2132),
.w133(w2133),
.w134(w2134),
.w135(w2135),
.w136(w2136),
.w137(w2137),
.w138(w2138),
.w139(w2139),
.w140(w2140),
.w141(w2141),
.w142(w2142),
.w143(w2143),
.w144(w2144),
.w145(w2145),
.w146(w2146),
.w147(w2147),
.w148(w2148),
.w20(w220),
.w21(w221),
.w22(w222),
.w23(w223),
.w24(w224),
.w25(w225),
.w26(w226),
.w27(w227),
.w28(w228),
.w29(w229),
.w210(w2210),
.w211(w2211),
.w212(w2212),
.w213(w2213),
.w214(w2214),
.w215(w2215),
.w216(w2216),
.w217(w2217),
.w218(w2218),
.w219(w2219),
.w220(w2220),
.w221(w2221),
.w222(w2222),
.w223(w2223),
.w224(w2224),
.w225(w2225),
.w226(w2226),
.w227(w2227),
.w228(w2228),
.w229(w2229),
.w230(w2230),
.w231(w2231),
.w232(w2232),
.w233(w2233),
.w234(w2234),
.w235(w2235),
.w236(w2236),
.w237(w2237),
.w238(w2238),
.w239(w2239),
.w240(w2240),
.w241(w2241),
.w242(w2242),
.w243(w2243),
.w244(w2244),
.w245(w2245),
.w246(w2246),
.w247(w2247),
.w248(w2248),
.bias(bias_2)
) block_1kernel_2
(
.clk(clk),
.rst(rst),
.valid_in(valid_in),
.In_0(In_0),
.In_1(In_1),
.In_2(In_2),
.Out(save_Out_2),
.valid_out(valid_out_2)
);

 
CONV_2D_1_Kernel_3_Channel_7 #(
.IMG_Width(IMG_Width), 
.IMG_Height(IMG_Height), 
.Datawidth(Datawidth), 
.Stride(Stride),
.ReLU(ReLU),
.w00(w300),
.w01(w301),
.w02(w302),
.w03(w303),
.w04(w304),
.w05(w305),
.w06(w306),
.w07(w307),
.w08(w308),
.w09(w309),
.w010(w3010),
.w011(w3011),
.w012(w3012),
.w013(w3013),
.w014(w3014),
.w015(w3015),
.w016(w3016),
.w017(w3017),
.w018(w3018),
.w019(w3019),
.w020(w3020),
.w021(w3021),
.w022(w3022),
.w023(w3023),
.w024(w3024),
.w025(w3025),
.w026(w3026),
.w027(w3027),
.w028(w3028),
.w029(w3029),
.w030(w3030),
.w031(w3031),
.w032(w3032),
.w033(w3033),
.w034(w3034),
.w035(w3035),
.w036(w3036),
.w037(w3037),
.w038(w3038),
.w039(w3039),
.w040(w3040),
.w041(w3041),
.w042(w3042),
.w043(w3043),
.w044(w3044),
.w045(w3045),
.w046(w3046),
.w047(w3047),
.w048(w3048),
.w10(w310),
.w11(w311),
.w12(w312),
.w13(w313),
.w14(w314),
.w15(w315),
.w16(w316),
.w17(w317),
.w18(w318),
.w19(w319),
.w110(w3110),
.w111(w3111),
.w112(w3112),
.w113(w3113),
.w114(w3114),
.w115(w3115),
.w116(w3116),
.w117(w3117),
.w118(w3118),
.w119(w3119),
.w120(w3120),
.w121(w3121),
.w122(w3122),
.w123(w3123),
.w124(w3124),
.w125(w3125),
.w126(w3126),
.w127(w3127),
.w128(w3128),
.w129(w3129),
.w130(w3130),
.w131(w3131),
.w132(w3132),
.w133(w3133),
.w134(w3134),
.w135(w3135),
.w136(w3136),
.w137(w3137),
.w138(w3138),
.w139(w3139),
.w140(w3140),
.w141(w3141),
.w142(w3142),
.w143(w3143),
.w144(w3144),
.w145(w3145),
.w146(w3146),
.w147(w3147),
.w148(w3148),
.w20(w320),
.w21(w321),
.w22(w322),
.w23(w323),
.w24(w324),
.w25(w325),
.w26(w326),
.w27(w327),
.w28(w328),
.w29(w329),
.w210(w3210),
.w211(w3211),
.w212(w3212),
.w213(w3213),
.w214(w3214),
.w215(w3215),
.w216(w3216),
.w217(w3217),
.w218(w3218),
.w219(w3219),
.w220(w3220),
.w221(w3221),
.w222(w3222),
.w223(w3223),
.w224(w3224),
.w225(w3225),
.w226(w3226),
.w227(w3227),
.w228(w3228),
.w229(w3229),
.w230(w3230),
.w231(w3231),
.w232(w3232),
.w233(w3233),
.w234(w3234),
.w235(w3235),
.w236(w3236),
.w237(w3237),
.w238(w3238),
.w239(w3239),
.w240(w3240),
.w241(w3241),
.w242(w3242),
.w243(w3243),
.w244(w3244),
.w245(w3245),
.w246(w3246),
.w247(w3247),
.w248(w3248),
.bias(bias_3)
) block_1kernel_3
(
.clk(clk),
.rst(rst),
.valid_in(valid_in),
.In_0(In_0),
.In_1(In_1),
.In_2(In_2),
.Out(save_Out_3),
.valid_out(valid_out_3)
);


endmodule 